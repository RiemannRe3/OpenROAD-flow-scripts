VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO SmallBuffer128
  FOREIGN SmallBuffer128 0 0 ;
  CLASS BLOCK ;
  SIZE 157.35 BY 188.415 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 162.7 115.38 164.1 ;
        RECT  2.9 122.7 115.38 124.1 ;
        RECT  2.9 82.7 115.38 84.1 ;
        RECT  2.9 42.7 115.38 44.1 ;
        RECT  2.9 2.7 115.38 4.1 ;
      LAYER metal4 ;
        RECT  114.9 1.315 115.38 186.285 ;
        RECT  58.9 1.315 59.38 186.285 ;
        RECT  2.9 1.315 3.38 186.285 ;
      LAYER metal1 ;
        RECT  1.14 186.115 156.18 186.285 ;
        RECT  1.14 183.315 156.18 183.485 ;
        RECT  1.14 180.515 156.18 180.685 ;
        RECT  1.14 177.715 156.18 177.885 ;
        RECT  1.14 174.915 156.18 175.085 ;
        RECT  1.14 172.115 156.18 172.285 ;
        RECT  1.14 169.315 156.18 169.485 ;
        RECT  1.14 166.515 156.18 166.685 ;
        RECT  1.14 163.715 156.18 163.885 ;
        RECT  1.14 160.915 156.18 161.085 ;
        RECT  1.14 158.115 156.18 158.285 ;
        RECT  1.14 155.315 156.18 155.485 ;
        RECT  1.14 152.515 156.18 152.685 ;
        RECT  1.14 149.715 156.18 149.885 ;
        RECT  1.14 146.915 156.18 147.085 ;
        RECT  1.14 144.115 156.18 144.285 ;
        RECT  1.14 141.315 156.18 141.485 ;
        RECT  1.14 138.515 156.18 138.685 ;
        RECT  1.14 135.715 156.18 135.885 ;
        RECT  1.14 132.915 156.18 133.085 ;
        RECT  1.14 130.115 156.18 130.285 ;
        RECT  1.14 127.315 156.18 127.485 ;
        RECT  1.14 124.515 156.18 124.685 ;
        RECT  1.14 121.715 156.18 121.885 ;
        RECT  1.14 118.915 156.18 119.085 ;
        RECT  1.14 116.115 156.18 116.285 ;
        RECT  1.14 113.315 156.18 113.485 ;
        RECT  1.14 110.515 156.18 110.685 ;
        RECT  1.14 107.715 156.18 107.885 ;
        RECT  1.14 104.915 156.18 105.085 ;
        RECT  1.14 102.115 156.18 102.285 ;
        RECT  1.14 99.315 156.18 99.485 ;
        RECT  1.14 96.515 156.18 96.685 ;
        RECT  1.14 93.715 156.18 93.885 ;
        RECT  1.14 90.915 156.18 91.085 ;
        RECT  1.14 88.115 156.18 88.285 ;
        RECT  1.14 85.315 156.18 85.485 ;
        RECT  1.14 82.515 156.18 82.685 ;
        RECT  1.14 79.715 156.18 79.885 ;
        RECT  1.14 76.915 156.18 77.085 ;
        RECT  1.14 74.115 156.18 74.285 ;
        RECT  1.14 71.315 156.18 71.485 ;
        RECT  1.14 68.515 156.18 68.685 ;
        RECT  1.14 65.715 156.18 65.885 ;
        RECT  1.14 62.915 156.18 63.085 ;
        RECT  1.14 60.115 156.18 60.285 ;
        RECT  1.14 57.315 156.18 57.485 ;
        RECT  1.14 54.515 156.18 54.685 ;
        RECT  1.14 51.715 156.18 51.885 ;
        RECT  1.14 48.915 156.18 49.085 ;
        RECT  1.14 46.115 156.18 46.285 ;
        RECT  1.14 43.315 156.18 43.485 ;
        RECT  1.14 40.515 156.18 40.685 ;
        RECT  1.14 37.715 156.18 37.885 ;
        RECT  1.14 34.915 156.18 35.085 ;
        RECT  1.14 32.115 156.18 32.285 ;
        RECT  1.14 29.315 156.18 29.485 ;
        RECT  1.14 26.515 156.18 26.685 ;
        RECT  1.14 23.715 156.18 23.885 ;
        RECT  1.14 20.915 156.18 21.085 ;
        RECT  1.14 18.115 156.18 18.285 ;
        RECT  1.14 15.315 156.18 15.485 ;
        RECT  1.14 12.515 156.18 12.685 ;
        RECT  1.14 9.715 156.18 9.885 ;
        RECT  1.14 6.915 156.18 7.085 ;
        RECT  1.14 4.115 156.18 4.285 ;
        RECT  1.14 1.315 156.18 1.485 ;
      VIA 115.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 186.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 186.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 186.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 183.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 183.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 183.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 180.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 180.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 180.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 177.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 177.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 177.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 175 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 175 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 175 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 172.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 172.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 172.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 186.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 186.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 186.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 183.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 183.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 183.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 180.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 180.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 180.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 177.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 177.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 177.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 175 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 175 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 175 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 172.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 172.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 172.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 186.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 186.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 186.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 183.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 183.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 183.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 180.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 180.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 180.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 177.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 177.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 177.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 175 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 175 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 175 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 172.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 172.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 172.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 182.7 143.38 184.1 ;
        RECT  30.9 142.7 143.38 144.1 ;
        RECT  30.9 102.7 143.38 104.1 ;
        RECT  30.9 62.7 143.38 64.1 ;
        RECT  30.9 22.7 143.38 24.1 ;
      LAYER metal4 ;
        RECT  142.9 2.715 143.38 184.885 ;
        RECT  86.9 2.715 87.38 184.885 ;
        RECT  30.9 2.715 31.38 184.885 ;
      LAYER metal1 ;
        RECT  1.14 184.715 156.18 184.885 ;
        RECT  1.14 181.915 156.18 182.085 ;
        RECT  1.14 179.115 156.18 179.285 ;
        RECT  1.14 176.315 156.18 176.485 ;
        RECT  1.14 173.515 156.18 173.685 ;
        RECT  1.14 170.715 156.18 170.885 ;
        RECT  1.14 167.915 156.18 168.085 ;
        RECT  1.14 165.115 156.18 165.285 ;
        RECT  1.14 162.315 156.18 162.485 ;
        RECT  1.14 159.515 156.18 159.685 ;
        RECT  1.14 156.715 156.18 156.885 ;
        RECT  1.14 153.915 156.18 154.085 ;
        RECT  1.14 151.115 156.18 151.285 ;
        RECT  1.14 148.315 156.18 148.485 ;
        RECT  1.14 145.515 156.18 145.685 ;
        RECT  1.14 142.715 156.18 142.885 ;
        RECT  1.14 139.915 156.18 140.085 ;
        RECT  1.14 137.115 156.18 137.285 ;
        RECT  1.14 134.315 156.18 134.485 ;
        RECT  1.14 131.515 156.18 131.685 ;
        RECT  1.14 128.715 156.18 128.885 ;
        RECT  1.14 125.915 156.18 126.085 ;
        RECT  1.14 123.115 156.18 123.285 ;
        RECT  1.14 120.315 156.18 120.485 ;
        RECT  1.14 117.515 156.18 117.685 ;
        RECT  1.14 114.715 156.18 114.885 ;
        RECT  1.14 111.915 156.18 112.085 ;
        RECT  1.14 109.115 156.18 109.285 ;
        RECT  1.14 106.315 156.18 106.485 ;
        RECT  1.14 103.515 156.18 103.685 ;
        RECT  1.14 100.715 156.18 100.885 ;
        RECT  1.14 97.915 156.18 98.085 ;
        RECT  1.14 95.115 156.18 95.285 ;
        RECT  1.14 92.315 156.18 92.485 ;
        RECT  1.14 89.515 156.18 89.685 ;
        RECT  1.14 86.715 156.18 86.885 ;
        RECT  1.14 83.915 156.18 84.085 ;
        RECT  1.14 81.115 156.18 81.285 ;
        RECT  1.14 78.315 156.18 78.485 ;
        RECT  1.14 75.515 156.18 75.685 ;
        RECT  1.14 72.715 156.18 72.885 ;
        RECT  1.14 69.915 156.18 70.085 ;
        RECT  1.14 67.115 156.18 67.285 ;
        RECT  1.14 64.315 156.18 64.485 ;
        RECT  1.14 61.515 156.18 61.685 ;
        RECT  1.14 58.715 156.18 58.885 ;
        RECT  1.14 55.915 156.18 56.085 ;
        RECT  1.14 53.115 156.18 53.285 ;
        RECT  1.14 50.315 156.18 50.485 ;
        RECT  1.14 47.515 156.18 47.685 ;
        RECT  1.14 44.715 156.18 44.885 ;
        RECT  1.14 41.915 156.18 42.085 ;
        RECT  1.14 39.115 156.18 39.285 ;
        RECT  1.14 36.315 156.18 36.485 ;
        RECT  1.14 33.515 156.18 33.685 ;
        RECT  1.14 30.715 156.18 30.885 ;
        RECT  1.14 27.915 156.18 28.085 ;
        RECT  1.14 25.115 156.18 25.285 ;
        RECT  1.14 22.315 156.18 22.485 ;
        RECT  1.14 19.515 156.18 19.685 ;
        RECT  1.14 16.715 156.18 16.885 ;
        RECT  1.14 13.915 156.18 14.085 ;
        RECT  1.14 11.115 156.18 11.285 ;
        RECT  1.14 8.315 156.18 8.485 ;
        RECT  1.14 5.515 156.18 5.685 ;
        RECT  1.14 2.715 156.18 2.885 ;
      VIA 143.14 183.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 183.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 183.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 183.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 183.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 183.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 183.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 183.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 183.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 184.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 184.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 184.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 182 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 182 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 182 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 179.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 179.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 179.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 176.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 176.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 176.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 173.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 173.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 173.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 170.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 170.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 170.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 184.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 184.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 184.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 182 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 182 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 182 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 179.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 179.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 179.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 176.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 176.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 176.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 173.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 173.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 173.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 170.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 170.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 170.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 184.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 184.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 184.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 182 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 182 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 182 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 179.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 179.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 179.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 176.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 176.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 176.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 173.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 173.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 173.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 170.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 170.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 170.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  31.945 0 32.085 0.14 ;
    END
  END clk
  PIN enable_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  157.21 53.76 157.35 53.9 ;
    END
  END enable_write
  PIN read_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  76.745 188.275 76.885 188.415 ;
    END
  END read_data[0]
  PIN read_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  76.185 0 76.325 0.14 ;
    END
  END read_data[1]
  PIN read_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  77.305 0 77.445 0.14 ;
    END
  END read_data[2]
  PIN read_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  83.465 188.275 83.605 188.415 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 98.56 0.14 98.7 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  77.865 0 78.005 0.14 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  82.905 188.275 83.045 188.415 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  80.665 188.275 80.805 188.415 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  82.345 188.275 82.485 188.415 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  75.625 0 75.765 0.14 ;
    END
  END read_data[9]
  PIN read_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  34.745 0 34.885 0.14 ;
    END
  END read_index[0]
  PIN read_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  122.105 188.275 122.245 188.415 ;
    END
  END read_index[1]
  PIN read_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  120.985 188.275 121.125 188.415 ;
    END
  END read_index[2]
  PIN read_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  120.425 188.275 120.565 188.415 ;
    END
  END read_index[3]
  PIN read_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  95.785 188.275 95.925 188.415 ;
    END
  END read_index[4]
  PIN read_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 128.8 0.14 128.94 ;
    END
  END read_index[5]
  PIN read_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 99.68 0.14 99.82 ;
    END
  END read_index[6]
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  77.305 188.275 77.445 188.415 ;
    END
  END write_data[0]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.225 188.275 81.365 188.415 ;
    END
  END write_data[1]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.425 188.275 78.565 188.415 ;
    END
  END write_data[2]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 132.16 0.14 132.3 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  71.705 188.275 71.845 188.415 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  79.545 188.275 79.685 188.415 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.985 188.275 79.125 188.415 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  80.105 188.275 80.245 188.415 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.785 188.275 81.925 188.415 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  77.865 188.275 78.005 188.415 ;
    END
  END write_data[9]
  PIN write_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  157.21 73.36 157.35 73.5 ;
    END
  END write_index[0]
  PIN write_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  157.21 72.24 157.35 72.38 ;
    END
  END write_index[1]
  PIN write_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  157.21 72.8 157.35 72.94 ;
    END
  END write_index[2]
  PIN write_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  72.825 0 72.965 0.14 ;
    END
  END write_index[3]
  PIN write_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  73.385 0 73.525 0.14 ;
    END
  END write_index[4]
  PIN write_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.425 0 78.565 0.14 ;
    END
  END write_index[5]
  PIN write_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.985 0 79.125 0.14 ;
    END
  END write_index[6]
  OBS
    LAYER metal1 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal2 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal3 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal4 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal5 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal6 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal7 ;
     RECT  0 0 157.35 188.415 ;
    LAYER metal8 ;
     RECT  0 0 157.35 188.415 ;
  END
END SmallBuffer128
END LIBRARY
