VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_960_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_960_340_1_3_300_300

VIA via2_3_960_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_960_340_1_3_320_320

VIA via3_4_960_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.045 0.035 ;
  ROWCOL 1 3 ;
END via3_4_960_340_1_3_320_320

VIA via4_5_960_2800_5_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0.02 0 0 0 ;
  ROWCOL 5 2 ;
END via4_5_960_2800_5_2_600_600

VIA via5_6_960_2800_5_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 5 2 ;
END via5_6_960_2800_5_2_600_600

VIA via6_7_960_2800_4_1_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.13 0.18 ;
  ROWCOL 4 1 ;
END via6_7_960_2800_4_1_600_600

MACRO myram
  FOREIGN myram 0 0 ;
  CLASS BLOCK ;
  SIZE 312.135 BY 157.07 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 152.7 283.38 154.1 ;
        RECT  2.9 122.7 283.38 124.1 ;
        RECT  2.9 92.7 283.38 94.1 ;
        RECT  2.9 62.7 283.38 64.1 ;
        RECT  2.9 32.7 283.38 34.1 ;
        RECT  2.9 2.7 283.38 4.1 ;
      LAYER metal4 ;
        RECT  282.9 1.315 283.38 155.485 ;
        RECT  226.9 1.315 227.38 155.485 ;
        RECT  170.9 1.315 171.38 155.485 ;
        RECT  114.9 1.315 115.38 155.485 ;
        RECT  58.9 1.315 59.38 155.485 ;
        RECT  2.9 1.315 3.38 155.485 ;
      LAYER metal1 ;
        RECT  1.14 155.315 311.03 155.485 ;
        RECT  1.14 152.515 311.03 152.685 ;
        RECT  1.14 149.715 311.03 149.885 ;
        RECT  1.14 146.915 311.03 147.085 ;
        RECT  1.14 144.115 311.03 144.285 ;
        RECT  1.14 141.315 311.03 141.485 ;
        RECT  1.14 138.515 311.03 138.685 ;
        RECT  1.14 135.715 311.03 135.885 ;
        RECT  1.14 132.915 311.03 133.085 ;
        RECT  1.14 130.115 311.03 130.285 ;
        RECT  1.14 127.315 311.03 127.485 ;
        RECT  1.14 124.515 311.03 124.685 ;
        RECT  1.14 121.715 311.03 121.885 ;
        RECT  1.14 118.915 311.03 119.085 ;
        RECT  1.14 116.115 311.03 116.285 ;
        RECT  1.14 113.315 311.03 113.485 ;
        RECT  1.14 110.515 311.03 110.685 ;
        RECT  1.14 107.715 311.03 107.885 ;
        RECT  1.14 104.915 311.03 105.085 ;
        RECT  1.14 102.115 311.03 102.285 ;
        RECT  1.14 99.315 311.03 99.485 ;
        RECT  1.14 96.515 311.03 96.685 ;
        RECT  1.14 93.715 311.03 93.885 ;
        RECT  1.14 90.915 311.03 91.085 ;
        RECT  1.14 88.115 311.03 88.285 ;
        RECT  1.14 85.315 311.03 85.485 ;
        RECT  1.14 82.515 311.03 82.685 ;
        RECT  1.14 79.715 311.03 79.885 ;
        RECT  1.14 76.915 311.03 77.085 ;
        RECT  1.14 74.115 311.03 74.285 ;
        RECT  1.14 71.315 311.03 71.485 ;
        RECT  1.14 68.515 311.03 68.685 ;
        RECT  1.14 65.715 311.03 65.885 ;
        RECT  1.14 62.915 311.03 63.085 ;
        RECT  1.14 60.115 311.03 60.285 ;
        RECT  1.14 57.315 311.03 57.485 ;
        RECT  1.14 54.515 311.03 54.685 ;
        RECT  1.14 51.715 311.03 51.885 ;
        RECT  1.14 48.915 311.03 49.085 ;
        RECT  1.14 46.115 311.03 46.285 ;
        RECT  1.14 43.315 311.03 43.485 ;
        RECT  1.14 40.515 311.03 40.685 ;
        RECT  1.14 37.715 311.03 37.885 ;
        RECT  1.14 34.915 311.03 35.085 ;
        RECT  1.14 32.115 311.03 32.285 ;
        RECT  1.14 29.315 311.03 29.485 ;
        RECT  1.14 26.515 311.03 26.685 ;
        RECT  1.14 23.715 311.03 23.885 ;
        RECT  1.14 20.915 311.03 21.085 ;
        RECT  1.14 18.115 311.03 18.285 ;
        RECT  1.14 15.315 311.03 15.485 ;
        RECT  1.14 12.515 311.03 12.685 ;
        RECT  1.14 9.715 311.03 9.885 ;
        RECT  1.14 6.915 311.03 7.085 ;
        RECT  1.14 4.115 311.03 4.285 ;
        RECT  1.14 1.315 311.03 1.485 ;
      VIA 283.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 153.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 153.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 153.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 93.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 93.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 93.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 137.7 255.38 139.1 ;
        RECT  30.9 107.7 255.38 109.1 ;
        RECT  30.9 77.7 255.38 79.1 ;
        RECT  30.9 47.7 255.38 49.1 ;
        RECT  30.9 17.7 255.38 19.1 ;
      LAYER metal4 ;
        RECT  254.9 2.715 255.38 154.085 ;
        RECT  198.9 2.715 199.38 154.085 ;
        RECT  142.9 2.715 143.38 154.085 ;
        RECT  86.9 2.715 87.38 154.085 ;
        RECT  30.9 2.715 31.38 154.085 ;
      LAYER metal1 ;
        RECT  1.14 153.915 311.03 154.085 ;
        RECT  1.14 151.115 311.03 151.285 ;
        RECT  1.14 148.315 311.03 148.485 ;
        RECT  1.14 145.515 311.03 145.685 ;
        RECT  1.14 142.715 311.03 142.885 ;
        RECT  1.14 139.915 311.03 140.085 ;
        RECT  1.14 137.115 311.03 137.285 ;
        RECT  1.14 134.315 311.03 134.485 ;
        RECT  1.14 131.515 311.03 131.685 ;
        RECT  1.14 128.715 311.03 128.885 ;
        RECT  1.14 125.915 311.03 126.085 ;
        RECT  1.14 123.115 311.03 123.285 ;
        RECT  1.14 120.315 311.03 120.485 ;
        RECT  1.14 117.515 311.03 117.685 ;
        RECT  1.14 114.715 311.03 114.885 ;
        RECT  1.14 111.915 311.03 112.085 ;
        RECT  1.14 109.115 311.03 109.285 ;
        RECT  1.14 106.315 311.03 106.485 ;
        RECT  1.14 103.515 311.03 103.685 ;
        RECT  1.14 100.715 311.03 100.885 ;
        RECT  1.14 97.915 311.03 98.085 ;
        RECT  1.14 95.115 311.03 95.285 ;
        RECT  1.14 92.315 311.03 92.485 ;
        RECT  1.14 89.515 311.03 89.685 ;
        RECT  1.14 86.715 311.03 86.885 ;
        RECT  1.14 83.915 311.03 84.085 ;
        RECT  1.14 81.115 311.03 81.285 ;
        RECT  1.14 78.315 311.03 78.485 ;
        RECT  1.14 75.515 311.03 75.685 ;
        RECT  1.14 72.715 311.03 72.885 ;
        RECT  1.14 69.915 311.03 70.085 ;
        RECT  1.14 67.115 311.03 67.285 ;
        RECT  1.14 64.315 311.03 64.485 ;
        RECT  1.14 61.515 311.03 61.685 ;
        RECT  1.14 58.715 311.03 58.885 ;
        RECT  1.14 55.915 311.03 56.085 ;
        RECT  1.14 53.115 311.03 53.285 ;
        RECT  1.14 50.315 311.03 50.485 ;
        RECT  1.14 47.515 311.03 47.685 ;
        RECT  1.14 44.715 311.03 44.885 ;
        RECT  1.14 41.915 311.03 42.085 ;
        RECT  1.14 39.115 311.03 39.285 ;
        RECT  1.14 36.315 311.03 36.485 ;
        RECT  1.14 33.515 311.03 33.685 ;
        RECT  1.14 30.715 311.03 30.885 ;
        RECT  1.14 27.915 311.03 28.085 ;
        RECT  1.14 25.115 311.03 25.285 ;
        RECT  1.14 22.315 311.03 22.485 ;
        RECT  1.14 19.515 311.03 19.685 ;
        RECT  1.14 16.715 311.03 16.885 ;
        RECT  1.14 13.915 311.03 14.085 ;
        RECT  1.14 11.115 311.03 11.285 ;
        RECT  1.14 8.315 311.03 8.485 ;
        RECT  1.14 5.515 311.03 5.685 ;
        RECT  1.14 2.715 311.03 2.885 ;
      VIA 255.14 138.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 138.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 138.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 108.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 108.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 108.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 78.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 78.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 78.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 138.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 138.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 138.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 108.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 108.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 108.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 78.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 78.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 78.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 138.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 138.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 138.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 108.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 108.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 108.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 78.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 78.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 78.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 138.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 138.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 138.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 108.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 108.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 108.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 78.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 78.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 78.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 138.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 138.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 138.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 108.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 108.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 108.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 78.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 78.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 78.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  161.305 156.93 161.445 157.07 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  2.825 156.93 2.965 157.07 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 6.16 312.135 6.3 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  301.305 0 301.445 0.14 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  285.625 0 285.765 0.14 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  190.425 0 190.565 0.14 ;
    END
  END addr_in[7]
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 117.04 312.135 117.18 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  208.905 156.93 209.045 157.07 ;
    END
  END clk
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 132.72 312.135 132.86 ;
    END
  END rd_out[0]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  253.705 0 253.845 0.14 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  97.465 156.93 97.605 157.07 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 69.44 312.135 69.58 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  34.185 156.93 34.325 157.07 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.105 156.93 66.245 157.07 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  192.665 156.93 192.805 157.07 ;
    END
  END rd_out[15]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  272.185 156.93 272.325 157.07 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  174.745 0 174.885 0.14 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 63.84 0.14 63.98 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  129.385 156.93 129.525 157.07 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 53.76 312.135 53.9 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  142.825 0 142.965 0.14 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  255.945 156.93 256.085 157.07 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  206.105 0 206.245 0.14 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  238.025 0 238.165 0.14 ;
    END
  END rd_out[9]
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  127.145 0 127.285 0.14 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  269.945 0 270.085 0.14 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  303.545 156.93 303.685 157.07 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  240.265 156.93 240.405 157.07 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  79.545 0 79.685 0.14 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.785 156.93 81.925 157.07 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  18.505 156.93 18.645 157.07 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 127.12 0.14 127.26 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 47.6 0.14 47.74 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 95.2 0.14 95.34 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  224.585 156.93 224.725 157.07 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 31.92 0.14 32.06 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 100.8 312.135 100.94 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 148.4 312.135 148.54 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  95.225 0 95.365 0.14 ;
    END
  END w_mask_in[9]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 85.12 312.135 85.26 ;
    END
  END wd_in[0]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  222.345 0 222.485 0.14 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  176.985 156.93 177.125 157.07 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 21.84 312.135 21.98 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  31.945 0 32.085 0.14 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  63.865 0 64.005 0.14 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 142.8 0.14 142.94 ;
    END
  END wd_in[15]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 16.24 0.14 16.38 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  111.465 0 111.605 0.14 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 111.44 0.14 111.58 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  287.865 156.93 288.005 157.07 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  113.705 156.93 113.845 157.07 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  145.065 156.93 145.205 157.07 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  159.065 0 159.205 0.14 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 79.52 0.14 79.66 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 156.93 50.005 157.07 ;
    END
  END wd_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  311.995 37.52 312.135 37.66 ;
    END
  END we_in
  OBS
    LAYER metal1 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal2 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal3 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal4 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal5 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal6 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal7 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal8 ;
     RECT  0 0 312.135 157.07 ;
    LAYER metal9 ;
     RECT  0 0 312.135 157.07 ;
  END
END myram
END LIBRARY
