VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_960_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_960_340_1_3_300_300

VIA via2_3_960_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_960_340_1_3_320_320

VIA via3_4_960_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.045 0.035 ;
  ROWCOL 1 3 ;
END via3_4_960_340_1_3_320_320

VIA via4_5_960_2800_5_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0.02 0 0 0 ;
  ROWCOL 5 2 ;
END via4_5_960_2800_5_2_600_600

VIA via5_6_960_2800_5_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 5 2 ;
END via5_6_960_2800_5_2_600_600

VIA via6_7_960_2800_4_1_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.13 0.18 ;
  ROWCOL 4 1 ;
END via6_7_960_2800_4_1_600_600

MACRO dctub_part1
  FOREIGN dctub_part1 0 0 ;
  CLASS BLOCK ;
  SIZE 143.485 BY 72.74 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 62.7 115.38 64.1 ;
        RECT  2.9 32.7 115.38 34.1 ;
        RECT  2.9 2.7 115.38 4.1 ;
      LAYER metal4 ;
        RECT  114.9 1.315 115.38 71.485 ;
        RECT  58.9 1.315 59.38 71.485 ;
        RECT  2.9 1.315 3.38 71.485 ;
      LAYER metal1 ;
        RECT  1.14 71.315 142.31 71.485 ;
        RECT  1.14 68.515 142.31 68.685 ;
        RECT  1.14 65.715 142.31 65.885 ;
        RECT  1.14 62.915 142.31 63.085 ;
        RECT  1.14 60.115 142.31 60.285 ;
        RECT  1.14 57.315 142.31 57.485 ;
        RECT  1.14 54.515 142.31 54.685 ;
        RECT  1.14 51.715 142.31 51.885 ;
        RECT  1.14 48.915 142.31 49.085 ;
        RECT  1.14 46.115 142.31 46.285 ;
        RECT  1.14 43.315 142.31 43.485 ;
        RECT  1.14 40.515 142.31 40.685 ;
        RECT  1.14 37.715 142.31 37.885 ;
        RECT  1.14 34.915 142.31 35.085 ;
        RECT  1.14 32.115 142.31 32.285 ;
        RECT  1.14 29.315 142.31 29.485 ;
        RECT  1.14 26.515 142.31 26.685 ;
        RECT  1.14 23.715 142.31 23.885 ;
        RECT  1.14 20.915 142.31 21.085 ;
        RECT  1.14 18.115 142.31 18.285 ;
        RECT  1.14 15.315 142.31 15.485 ;
        RECT  1.14 12.515 142.31 12.685 ;
        RECT  1.14 9.715 142.31 9.885 ;
        RECT  1.14 6.915 142.31 7.085 ;
        RECT  1.14 4.115 142.31 4.285 ;
        RECT  1.14 1.315 142.31 1.485 ;
      VIA 115.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 47.7 87.38 49.1 ;
        RECT  30.9 17.7 87.38 19.1 ;
      LAYER metal4 ;
        RECT  86.9 2.715 87.38 70.085 ;
        RECT  30.9 2.715 31.38 70.085 ;
      LAYER metal1 ;
        RECT  1.14 69.915 142.31 70.085 ;
        RECT  1.14 67.115 142.31 67.285 ;
        RECT  1.14 64.315 142.31 64.485 ;
        RECT  1.14 61.515 142.31 61.685 ;
        RECT  1.14 58.715 142.31 58.885 ;
        RECT  1.14 55.915 142.31 56.085 ;
        RECT  1.14 53.115 142.31 53.285 ;
        RECT  1.14 50.315 142.31 50.485 ;
        RECT  1.14 47.515 142.31 47.685 ;
        RECT  1.14 44.715 142.31 44.885 ;
        RECT  1.14 41.915 142.31 42.085 ;
        RECT  1.14 39.115 142.31 39.285 ;
        RECT  1.14 36.315 142.31 36.485 ;
        RECT  1.14 33.515 142.31 33.685 ;
        RECT  1.14 30.715 142.31 30.885 ;
        RECT  1.14 27.915 142.31 28.085 ;
        RECT  1.14 25.115 142.31 25.285 ;
        RECT  1.14 22.315 142.31 22.485 ;
        RECT  1.14 19.515 142.31 19.685 ;
        RECT  1.14 16.715 142.31 16.885 ;
        RECT  1.14 13.915 142.31 14.085 ;
        RECT  1.14 11.115 142.31 11.285 ;
        RECT  1.14 8.315 142.31 8.485 ;
        RECT  1.14 5.515 142.31 5.685 ;
        RECT  1.14 2.715 142.31 2.885 ;
      VIA 87.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  24.665 0 24.805 0.14 ;
    END
  END clk
  PIN ddgo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 64.96 0.14 65.1 ;
    END
  END ddgo
  PIN ddin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  89.065 0 89.205 0.14 ;
    END
  END ddin[1]
  PIN ddin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  41.465 72.6 41.605 72.74 ;
    END
  END ddin[2]
  PIN ddin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 19.6 143.485 19.74 ;
    END
  END ddin[3]
  PIN ddin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.225 0 81.365 0.14 ;
    END
  END ddin[4]
  PIN ddin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END ddin[5]
  PIN ddin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  9.545 72.6 9.685 72.74 ;
    END
  END ddin[6]
  PIN ddin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  33.625 72.6 33.765 72.74 ;
    END
  END ddin[7]
  PIN ddin[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  121.545 0 121.685 0.14 ;
    END
  END ddin[8]
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  106.425 72.6 106.565 72.74 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  113.145 0 113.285 0.14 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  122.105 72.6 122.245 72.74 ;
    END
  END dout0[11]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  129.385 0 129.525 0.14 ;
    END
  END dout0[1]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 72.6 50.005 72.74 ;
    END
  END dout0[2]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  137.785 0 137.925 0.14 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  1.145 72.6 1.285 72.74 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 59.92 143.485 60.06 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 32.48 0.14 32.62 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 48.72 0.14 48.86 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  17.385 72.6 17.525 72.74 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  105.305 0 105.445 0.14 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 56.56 0.14 56.7 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 43.68 143.485 43.82 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 16.24 0.14 16.38 ;
    END
  END dout1[11]
  PIN dout1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  98.025 72.6 98.165 72.74 ;
    END
  END dout1[1]
  PIN dout1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 24.64 0.14 24.78 ;
    END
  END dout1[2]
  PIN dout1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 67.76 143.485 67.9 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.785 72.6 81.925 72.74 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 27.44 143.485 27.58 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  114.265 72.6 114.405 72.74 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  8.425 0 8.565 0.14 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.105 72.6 66.245 72.74 ;
    END
  END dout1[9]
  PIN dout2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 51.52 143.485 51.66 ;
    END
  END dout2[0]
  PIN dout2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  40.905 0 41.045 0.14 ;
    END
  END dout2[10]
  PIN dout2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 35.84 143.485 35.98 ;
    END
  END dout2[11]
  PIN dout2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  96.905 0 97.045 0.14 ;
    END
  END dout2[1]
  PIN dout2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  90.185 72.6 90.325 72.74 ;
    END
  END dout2[2]
  PIN dout2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 3.36 143.485 3.5 ;
    END
  END dout2[3]
  PIN dout2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END dout2[4]
  PIN dout2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END dout2[5]
  PIN dout2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END dout2[6]
  PIN dout2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 8.4 0.14 8.54 ;
    END
  END dout2[7]
  PIN dout2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END dout2[8]
  PIN dout2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  138.345 72.6 138.485 72.74 ;
    END
  END dout2[9]
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  130.505 72.6 130.645 72.74 ;
    END
  END ena
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  57.705 72.6 57.845 72.74 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  73.945 72.6 74.085 72.74 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  72.825 0 72.965 0.14 ;
    END
  END x[2]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 40.88 0.14 41.02 ;
    END
  END y[0]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  25.225 72.6 25.365 72.74 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  143.345 11.2 143.485 11.34 ;
    END
  END y[2]
  OBS
    LAYER metal1 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal2 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal3 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal4 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal5 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal6 ;
     RECT  0 0 143.485 72.74 ;
    LAYER metal7 ;
     RECT  0 0 143.485 72.74 ;
  END
END dctub_part1
END LIBRARY
