VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_960_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_960_340_1_3_300_300

VIA via2_3_960_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_960_340_1_3_320_320

VIA via3_4_960_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.045 0.035 ;
  ROWCOL 1 3 ;
END via3_4_960_340_1_3_320_320

VIA via4_5_960_2800_5_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0.02 0 0 0 ;
  ROWCOL 5 2 ;
END via4_5_960_2800_5_2_600_600

VIA via5_6_960_2800_5_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 5 2 ;
END via5_6_960_2800_5_2_600_600

VIA via6_7_960_2800_4_1_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.13 0.18 ;
  ROWCOL 4 1 ;
END via6_7_960_2800_4_1_600_600

MACRO dctub_part3
  FOREIGN dctub_part3 0 0 ;
  CLASS BLOCK ;
  SIZE 98.66 BY 79.33 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 62.7 59.38 64.1 ;
        RECT  2.9 32.7 59.38 34.1 ;
        RECT  2.9 2.7 59.38 4.1 ;
      LAYER metal4 ;
        RECT  58.9 1.315 59.38 77.085 ;
        RECT  2.9 1.315 3.38 77.085 ;
      LAYER metal1 ;
        RECT  1.14 76.915 97.66 77.085 ;
        RECT  1.14 74.115 97.66 74.285 ;
        RECT  1.14 71.315 97.66 71.485 ;
        RECT  1.14 68.515 97.66 68.685 ;
        RECT  1.14 65.715 97.66 65.885 ;
        RECT  1.14 62.915 97.66 63.085 ;
        RECT  1.14 60.115 97.66 60.285 ;
        RECT  1.14 57.315 97.66 57.485 ;
        RECT  1.14 54.515 97.66 54.685 ;
        RECT  1.14 51.715 97.66 51.885 ;
        RECT  1.14 48.915 97.66 49.085 ;
        RECT  1.14 46.115 97.66 46.285 ;
        RECT  1.14 43.315 97.66 43.485 ;
        RECT  1.14 40.515 97.66 40.685 ;
        RECT  1.14 37.715 97.66 37.885 ;
        RECT  1.14 34.915 97.66 35.085 ;
        RECT  1.14 32.115 97.66 32.285 ;
        RECT  1.14 29.315 97.66 29.485 ;
        RECT  1.14 26.515 97.66 26.685 ;
        RECT  1.14 23.715 97.66 23.885 ;
        RECT  1.14 20.915 97.66 21.085 ;
        RECT  1.14 18.115 97.66 18.285 ;
        RECT  1.14 15.315 97.66 15.485 ;
        RECT  1.14 12.515 97.66 12.685 ;
        RECT  1.14 9.715 97.66 9.885 ;
        RECT  1.14 6.915 97.66 7.085 ;
        RECT  1.14 4.115 97.66 4.285 ;
        RECT  1.14 1.315 97.66 1.485 ;
      VIA 59.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 33.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 33.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 47.7 87.38 49.1 ;
        RECT  30.9 17.7 87.38 19.1 ;
      LAYER metal4 ;
        RECT  86.9 2.715 87.38 75.685 ;
        RECT  30.9 2.715 31.38 75.685 ;
      LAYER metal1 ;
        RECT  1.14 75.515 97.66 75.685 ;
        RECT  1.14 72.715 97.66 72.885 ;
        RECT  1.14 69.915 97.66 70.085 ;
        RECT  1.14 67.115 97.66 67.285 ;
        RECT  1.14 64.315 97.66 64.485 ;
        RECT  1.14 61.515 97.66 61.685 ;
        RECT  1.14 58.715 97.66 58.885 ;
        RECT  1.14 55.915 97.66 56.085 ;
        RECT  1.14 53.115 97.66 53.285 ;
        RECT  1.14 50.315 97.66 50.485 ;
        RECT  1.14 47.515 97.66 47.685 ;
        RECT  1.14 44.715 97.66 44.885 ;
        RECT  1.14 41.915 97.66 42.085 ;
        RECT  1.14 39.115 97.66 39.285 ;
        RECT  1.14 36.315 97.66 36.485 ;
        RECT  1.14 33.515 97.66 33.685 ;
        RECT  1.14 30.715 97.66 30.885 ;
        RECT  1.14 27.915 97.66 28.085 ;
        RECT  1.14 25.115 97.66 25.285 ;
        RECT  1.14 22.315 97.66 22.485 ;
        RECT  1.14 19.515 97.66 19.685 ;
        RECT  1.14 16.715 97.66 16.885 ;
        RECT  1.14 13.915 97.66 14.085 ;
        RECT  1.14 11.115 97.66 11.285 ;
        RECT  1.14 8.315 97.66 8.485 ;
        RECT  1.14 5.515 97.66 5.685 ;
        RECT  1.14 2.715 97.66 2.885 ;
      VIA 87.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 48.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 48.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 18.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 18.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  20.185 0 20.325 0.14 ;
    END
  END clk
  PIN ddgo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 53.2 0.14 53.34 ;
    END
  END ddgo
  PIN ddin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  73.385 0 73.525 0.14 ;
    END
  END ddin[1]
  PIN ddin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  14.585 79.19 14.725 79.33 ;
    END
  END ddin[2]
  PIN ddin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 35.28 98.66 35.42 ;
    END
  END ddin[3]
  PIN ddin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END ddin[4]
  PIN ddin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  53.225 0 53.365 0.14 ;
    END
  END ddin[5]
  PIN ddin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 66.64 0.14 66.78 ;
    END
  END ddin[6]
  PIN ddin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  8.425 79.19 8.565 79.33 ;
    END
  END ddin[7]
  PIN ddin[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 2.24 98.66 2.38 ;
    END
  END ddin[8]
  PIN dout5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  67.785 79.19 67.925 79.33 ;
    END
  END dout5[0]
  PIN dout5[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  92.985 0 93.125 0.14 ;
    END
  END dout5[10]
  PIN dout5[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  81.225 79.19 81.365 79.33 ;
    END
  END dout5[11]
  PIN dout5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 8.96 98.66 9.1 ;
    END
  END dout5[1]
  PIN dout5[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  21.305 79.19 21.445 79.33 ;
    END
  END dout5[2]
  PIN dout5[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 15.68 98.66 15.82 ;
    END
  END dout5[3]
  PIN dout5[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 59.92 0.14 60.06 ;
    END
  END dout5[4]
  PIN dout5[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 68.88 98.66 69.02 ;
    END
  END dout5[5]
  PIN dout5[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 26.88 0.14 27.02 ;
    END
  END dout5[6]
  PIN dout5[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 40.32 0.14 40.46 ;
    END
  END dout5[7]
  PIN dout5[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 73.36 0.14 73.5 ;
    END
  END dout5[8]
  PIN dout5[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  86.825 0 86.965 0.14 ;
    END
  END dout5[9]
  PIN dout6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 46.48 0.14 46.62 ;
    END
  END dout6[0]
  PIN dout6[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 55.44 98.66 55.58 ;
    END
  END dout6[10]
  PIN dout6[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 13.44 0.14 13.58 ;
    END
  END dout6[11]
  PIN dout6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  61.065 79.19 61.205 79.33 ;
    END
  END dout6[1]
  PIN dout6[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 20.16 0.14 20.3 ;
    END
  END dout6[2]
  PIN dout6[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 75.6 98.66 75.74 ;
    END
  END dout6[3]
  PIN dout6[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.185 79.19 48.325 79.33 ;
    END
  END dout6[4]
  PIN dout6[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 42 98.66 42.14 ;
    END
  END dout6[5]
  PIN dout6[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  74.505 79.19 74.645 79.33 ;
    END
  END dout6[6]
  PIN dout6[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  6.745 0 6.885 0.14 ;
    END
  END dout6[7]
  PIN dout6[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END dout6[8]
  PIN dout6[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  34.745 79.19 34.885 79.33 ;
    END
  END dout6[9]
  PIN dout7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 62.16 98.66 62.3 ;
    END
  END dout7[0]
  PIN dout7[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  33.625 0 33.765 0.14 ;
    END
  END dout7[10]
  PIN dout7[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 48.72 98.66 48.86 ;
    END
  END dout7[11]
  PIN dout7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  80.105 0 80.245 0.14 ;
    END
  END dout7[1]
  PIN dout7[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  54.345 79.19 54.485 79.33 ;
    END
  END dout7[2]
  PIN dout7[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 22.4 98.66 22.54 ;
    END
  END dout7[3]
  PIN dout7[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  13.465 0 13.605 0.14 ;
    END
  END dout7[4]
  PIN dout7[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.905 0 27.045 0.14 ;
    END
  END dout7[5]
  PIN dout7[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  40.345 0 40.485 0.14 ;
    END
  END dout7[6]
  PIN dout7[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 6.72 0.14 6.86 ;
    END
  END dout7[7]
  PIN dout7[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  46.505 0 46.645 0.14 ;
    END
  END dout7[8]
  PIN dout7[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  94.665 79.19 94.805 79.33 ;
    END
  END dout7[9]
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  87.945 79.19 88.085 79.33 ;
    END
  END ena
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  28.025 79.19 28.165 79.33 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  41.465 79.19 41.605 79.33 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END x[2]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 33.6 0.14 33.74 ;
    END
  END y[0]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  1.705 79.19 1.845 79.33 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  98.52 29.12 98.66 29.26 ;
    END
  END y[2]
  OBS
    LAYER metal1 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal2 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal3 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal4 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal5 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal6 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal7 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal8 ;
     RECT  0 0 98.66 79.33 ;
    LAYER metal9 ;
     RECT  0 0 98.66 79.33 ;
  END
END dctub_part3
END LIBRARY
