VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO SmallBuffer256
  FOREIGN SmallBuffer256 0 0 ;
  CLASS BLOCK ;
  SIZE 340.1 BY 171.615 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 162.7 339.38 164.1 ;
        RECT  2.9 122.7 339.38 124.1 ;
        RECT  2.9 82.7 339.38 84.1 ;
        RECT  2.9 42.7 339.38 44.1 ;
        RECT  2.9 2.7 339.38 4.1 ;
      LAYER metal4 ;
        RECT  338.9 1.315 339.38 169.485 ;
        RECT  282.9 1.315 283.38 169.485 ;
        RECT  226.9 1.315 227.38 169.485 ;
        RECT  170.9 1.315 171.38 169.485 ;
        RECT  114.9 1.315 115.38 169.485 ;
        RECT  58.9 1.315 59.38 169.485 ;
        RECT  2.9 1.315 3.38 169.485 ;
      LAYER metal1 ;
        RECT  1.14 169.315 340.1 169.485 ;
        RECT  1.14 166.515 340.1 166.685 ;
        RECT  1.14 163.715 340.1 163.885 ;
        RECT  1.14 160.915 340.1 161.085 ;
        RECT  1.14 158.115 340.1 158.285 ;
        RECT  1.14 155.315 340.1 155.485 ;
        RECT  1.14 152.515 340.1 152.685 ;
        RECT  1.14 149.715 340.1 149.885 ;
        RECT  1.14 146.915 340.1 147.085 ;
        RECT  1.14 144.115 340.1 144.285 ;
        RECT  1.14 141.315 340.1 141.485 ;
        RECT  1.14 138.515 340.1 138.685 ;
        RECT  1.14 135.715 340.1 135.885 ;
        RECT  1.14 132.915 340.1 133.085 ;
        RECT  1.14 130.115 340.1 130.285 ;
        RECT  1.14 127.315 340.1 127.485 ;
        RECT  1.14 124.515 340.1 124.685 ;
        RECT  1.14 121.715 340.1 121.885 ;
        RECT  1.14 118.915 340.1 119.085 ;
        RECT  1.14 116.115 340.1 116.285 ;
        RECT  1.14 113.315 340.1 113.485 ;
        RECT  1.14 110.515 340.1 110.685 ;
        RECT  1.14 107.715 340.1 107.885 ;
        RECT  1.14 104.915 340.1 105.085 ;
        RECT  1.14 102.115 340.1 102.285 ;
        RECT  1.14 99.315 340.1 99.485 ;
        RECT  1.14 96.515 340.1 96.685 ;
        RECT  1.14 93.715 340.1 93.885 ;
        RECT  1.14 90.915 340.1 91.085 ;
        RECT  1.14 88.115 340.1 88.285 ;
        RECT  1.14 85.315 340.1 85.485 ;
        RECT  1.14 82.515 340.1 82.685 ;
        RECT  1.14 79.715 340.1 79.885 ;
        RECT  1.14 76.915 340.1 77.085 ;
        RECT  1.14 74.115 340.1 74.285 ;
        RECT  1.14 71.315 340.1 71.485 ;
        RECT  1.14 68.515 340.1 68.685 ;
        RECT  1.14 65.715 340.1 65.885 ;
        RECT  1.14 62.915 340.1 63.085 ;
        RECT  1.14 60.115 340.1 60.285 ;
        RECT  1.14 57.315 340.1 57.485 ;
        RECT  1.14 54.515 340.1 54.685 ;
        RECT  1.14 51.715 340.1 51.885 ;
        RECT  1.14 48.915 340.1 49.085 ;
        RECT  1.14 46.115 340.1 46.285 ;
        RECT  1.14 43.315 340.1 43.485 ;
        RECT  1.14 40.515 340.1 40.685 ;
        RECT  1.14 37.715 340.1 37.885 ;
        RECT  1.14 34.915 340.1 35.085 ;
        RECT  1.14 32.115 340.1 32.285 ;
        RECT  1.14 29.315 340.1 29.485 ;
        RECT  1.14 26.515 340.1 26.685 ;
        RECT  1.14 23.715 340.1 23.885 ;
        RECT  1.14 20.915 340.1 21.085 ;
        RECT  1.14 18.115 340.1 18.285 ;
        RECT  1.14 15.315 340.1 15.485 ;
        RECT  1.14 12.515 340.1 12.685 ;
        RECT  1.14 9.715 340.1 9.885 ;
        RECT  1.14 6.915 340.1 7.085 ;
        RECT  1.14 4.115 340.1 4.285 ;
        RECT  1.14 1.315 340.1 1.485 ;
      VIA 339.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 339.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 339.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 339.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 339.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 339.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 339.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 339.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 339.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 339.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 339.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 339.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 339.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 339.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 339.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 283.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 283.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 283.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 227.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 227.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 227.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 171.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 171.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 171.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 115.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 339.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 339.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 339.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 339.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 283.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 283.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 283.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 227.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 227.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 227.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 171.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 171.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 171.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 115.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 115.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 142.7 311.38 144.1 ;
        RECT  30.9 102.7 311.38 104.1 ;
        RECT  30.9 62.7 311.38 64.1 ;
        RECT  30.9 22.7 311.38 24.1 ;
      LAYER metal4 ;
        RECT  310.9 2.715 311.38 168.085 ;
        RECT  254.9 2.715 255.38 168.085 ;
        RECT  198.9 2.715 199.38 168.085 ;
        RECT  142.9 2.715 143.38 168.085 ;
        RECT  86.9 2.715 87.38 168.085 ;
        RECT  30.9 2.715 31.38 168.085 ;
      LAYER metal1 ;
        RECT  1.14 167.915 340.1 168.085 ;
        RECT  1.14 165.115 340.1 165.285 ;
        RECT  1.14 162.315 340.1 162.485 ;
        RECT  1.14 159.515 340.1 159.685 ;
        RECT  1.14 156.715 340.1 156.885 ;
        RECT  1.14 153.915 340.1 154.085 ;
        RECT  1.14 151.115 340.1 151.285 ;
        RECT  1.14 148.315 340.1 148.485 ;
        RECT  1.14 145.515 340.1 145.685 ;
        RECT  1.14 142.715 340.1 142.885 ;
        RECT  1.14 139.915 340.1 140.085 ;
        RECT  1.14 137.115 340.1 137.285 ;
        RECT  1.14 134.315 340.1 134.485 ;
        RECT  1.14 131.515 340.1 131.685 ;
        RECT  1.14 128.715 340.1 128.885 ;
        RECT  1.14 125.915 340.1 126.085 ;
        RECT  1.14 123.115 340.1 123.285 ;
        RECT  1.14 120.315 340.1 120.485 ;
        RECT  1.14 117.515 340.1 117.685 ;
        RECT  1.14 114.715 340.1 114.885 ;
        RECT  1.14 111.915 340.1 112.085 ;
        RECT  1.14 109.115 340.1 109.285 ;
        RECT  1.14 106.315 340.1 106.485 ;
        RECT  1.14 103.515 340.1 103.685 ;
        RECT  1.14 100.715 340.1 100.885 ;
        RECT  1.14 97.915 340.1 98.085 ;
        RECT  1.14 95.115 340.1 95.285 ;
        RECT  1.14 92.315 340.1 92.485 ;
        RECT  1.14 89.515 340.1 89.685 ;
        RECT  1.14 86.715 340.1 86.885 ;
        RECT  1.14 83.915 340.1 84.085 ;
        RECT  1.14 81.115 340.1 81.285 ;
        RECT  1.14 78.315 340.1 78.485 ;
        RECT  1.14 75.515 340.1 75.685 ;
        RECT  1.14 72.715 340.1 72.885 ;
        RECT  1.14 69.915 340.1 70.085 ;
        RECT  1.14 67.115 340.1 67.285 ;
        RECT  1.14 64.315 340.1 64.485 ;
        RECT  1.14 61.515 340.1 61.685 ;
        RECT  1.14 58.715 340.1 58.885 ;
        RECT  1.14 55.915 340.1 56.085 ;
        RECT  1.14 53.115 340.1 53.285 ;
        RECT  1.14 50.315 340.1 50.485 ;
        RECT  1.14 47.515 340.1 47.685 ;
        RECT  1.14 44.715 340.1 44.885 ;
        RECT  1.14 41.915 340.1 42.085 ;
        RECT  1.14 39.115 340.1 39.285 ;
        RECT  1.14 36.315 340.1 36.485 ;
        RECT  1.14 33.515 340.1 33.685 ;
        RECT  1.14 30.715 340.1 30.885 ;
        RECT  1.14 27.915 340.1 28.085 ;
        RECT  1.14 25.115 340.1 25.285 ;
        RECT  1.14 22.315 340.1 22.485 ;
        RECT  1.14 19.515 340.1 19.685 ;
        RECT  1.14 16.715 340.1 16.885 ;
        RECT  1.14 13.915 340.1 14.085 ;
        RECT  1.14 11.115 340.1 11.285 ;
        RECT  1.14 8.315 340.1 8.485 ;
        RECT  1.14 5.515 340.1 5.685 ;
        RECT  1.14 2.715 340.1 2.885 ;
      VIA 311.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 311.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 311.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 311.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 311.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 311.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 311.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 311.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 311.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 311.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 311.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 311.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 255.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 255.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 255.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 199.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 199.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 199.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 143.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 143.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 143.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 143.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 143.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 103.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 103.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 311.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 311.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 311.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 311.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 255.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 255.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 255.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 199.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 199.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 199.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 143.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 143.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  228.505 171.475 228.645 171.615 ;
    END
  END clk
  PIN enable_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  164.105 171.475 164.245 171.615 ;
    END
  END enable_write
  PIN read_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  176.985 171.475 177.125 171.615 ;
    END
  END read_data[0]
  PIN read_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  183.145 171.475 183.285 171.615 ;
    END
  END read_data[1]
  PIN read_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  175.865 171.475 176.005 171.615 ;
    END
  END read_data[2]
  PIN read_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  185.945 171.475 186.085 171.615 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  174.745 171.475 174.885 171.615 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  185.385 171.475 185.525 171.615 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  182.585 171.475 182.725 171.615 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  180.345 171.475 180.485 171.615 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  175.305 171.475 175.445 171.615 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  174.185 171.475 174.325 171.615 ;
    END
  END read_data[9]
  PIN read_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  227.945 171.475 228.085 171.615 ;
    END
  END read_index[0]
  PIN read_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  227.385 171.475 227.525 171.615 ;
    END
  END read_index[1]
  PIN read_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  226.825 171.475 226.965 171.615 ;
    END
  END read_index[2]
  PIN read_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  226.265 171.475 226.405 171.615 ;
    END
  END read_index[3]
  PIN read_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  225.705 171.475 225.845 171.615 ;
    END
  END read_index[4]
  PIN read_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  112.585 0 112.725 0.14 ;
    END
  END read_index[5]
  PIN read_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  171.385 171.475 171.525 171.615 ;
    END
  END read_index[6]
  PIN read_index[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  182.025 171.475 182.165 171.615 ;
    END
  END read_index[7]
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  124.905 171.475 125.045 171.615 ;
    END
  END write_data[0]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  129.385 171.475 129.525 171.615 ;
    END
  END write_data[1]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  127.145 171.475 127.285 171.615 ;
    END
  END write_data[2]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  126.025 171.475 126.165 171.615 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  124.345 171.475 124.485 171.615 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  128.265 171.475 128.405 171.615 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  127.705 171.475 127.845 171.615 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  125.465 171.475 125.605 171.615 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  128.825 171.475 128.965 171.615 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  126.585 171.475 126.725 171.615 ;
    END
  END write_data[9]
  PIN write_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  116.505 0 116.645 0.14 ;
    END
  END write_index[0]
  PIN write_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  118.185 0 118.325 0.14 ;
    END
  END write_index[1]
  PIN write_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  117.065 0 117.205 0.14 ;
    END
  END write_index[2]
  PIN write_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  117.625 0 117.765 0.14 ;
    END
  END write_index[3]
  PIN write_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  165.225 171.475 165.365 171.615 ;
    END
  END write_index[4]
  PIN write_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  164.665 171.475 164.805 171.615 ;
    END
  END write_index[5]
  PIN write_index[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  162.985 171.475 163.125 171.615 ;
    END
  END write_index[6]
  PIN write_index[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  163.545 171.475 163.685 171.615 ;
    END
  END write_index[7]
  OBS
    LAYER metal1 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal2 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal3 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal4 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal5 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal6 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal7 ;
     RECT  1.14 0 340.1 171.615 ;
    LAYER metal9 ;
     RECT  1.14 0 340.1 171.615 ;
  END
END SmallBuffer256
END LIBRARY
