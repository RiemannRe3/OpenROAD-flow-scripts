VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO SmallBuffer64
  FOREIGN SmallBuffer64 0 0 ;
  CLASS BLOCK ;
  SIZE 71.785 BY 210.085 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 202.7 59.38 204.1 ;
        RECT  2.9 162.7 59.38 164.1 ;
        RECT  2.9 122.7 59.38 124.1 ;
        RECT  2.9 82.7 59.38 84.1 ;
        RECT  2.9 42.7 59.38 44.1 ;
        RECT  2.9 2.7 59.38 4.1 ;
      LAYER metal4 ;
        RECT  58.9 1.315 59.38 208.685 ;
        RECT  2.9 1.315 3.38 208.685 ;
      LAYER metal1 ;
        RECT  1.14 208.515 70.68 208.685 ;
        RECT  1.14 205.715 70.68 205.885 ;
        RECT  1.14 202.915 70.68 203.085 ;
        RECT  1.14 200.115 70.68 200.285 ;
        RECT  1.14 197.315 70.68 197.485 ;
        RECT  1.14 194.515 70.68 194.685 ;
        RECT  1.14 191.715 70.68 191.885 ;
        RECT  1.14 188.915 70.68 189.085 ;
        RECT  1.14 186.115 70.68 186.285 ;
        RECT  1.14 183.315 70.68 183.485 ;
        RECT  1.14 180.515 70.68 180.685 ;
        RECT  1.14 177.715 70.68 177.885 ;
        RECT  1.14 174.915 70.68 175.085 ;
        RECT  1.14 172.115 70.68 172.285 ;
        RECT  1.14 169.315 70.68 169.485 ;
        RECT  1.14 166.515 70.68 166.685 ;
        RECT  1.14 163.715 70.68 163.885 ;
        RECT  1.14 160.915 70.68 161.085 ;
        RECT  1.14 158.115 70.68 158.285 ;
        RECT  1.14 155.315 70.68 155.485 ;
        RECT  1.14 152.515 70.68 152.685 ;
        RECT  1.14 149.715 70.68 149.885 ;
        RECT  1.14 146.915 70.68 147.085 ;
        RECT  1.14 144.115 70.68 144.285 ;
        RECT  1.14 141.315 70.68 141.485 ;
        RECT  1.14 138.515 70.68 138.685 ;
        RECT  1.14 135.715 70.68 135.885 ;
        RECT  1.14 132.915 70.68 133.085 ;
        RECT  1.14 130.115 70.68 130.285 ;
        RECT  1.14 127.315 70.68 127.485 ;
        RECT  1.14 124.515 70.68 124.685 ;
        RECT  1.14 121.715 70.68 121.885 ;
        RECT  1.14 118.915 70.68 119.085 ;
        RECT  1.14 116.115 70.68 116.285 ;
        RECT  1.14 113.315 70.68 113.485 ;
        RECT  1.14 110.515 70.68 110.685 ;
        RECT  1.14 107.715 70.68 107.885 ;
        RECT  1.14 104.915 70.68 105.085 ;
        RECT  1.14 102.115 70.68 102.285 ;
        RECT  1.14 99.315 70.68 99.485 ;
        RECT  1.14 96.515 70.68 96.685 ;
        RECT  1.14 93.715 70.68 93.885 ;
        RECT  1.14 90.915 70.68 91.085 ;
        RECT  1.14 88.115 70.68 88.285 ;
        RECT  1.14 85.315 70.68 85.485 ;
        RECT  1.14 82.515 70.68 82.685 ;
        RECT  1.14 79.715 70.68 79.885 ;
        RECT  1.14 76.915 70.68 77.085 ;
        RECT  1.14 74.115 70.68 74.285 ;
        RECT  1.14 71.315 70.68 71.485 ;
        RECT  1.14 68.515 70.68 68.685 ;
        RECT  1.14 65.715 70.68 65.885 ;
        RECT  1.14 62.915 70.68 63.085 ;
        RECT  1.14 60.115 70.68 60.285 ;
        RECT  1.14 57.315 70.68 57.485 ;
        RECT  1.14 54.515 70.68 54.685 ;
        RECT  1.14 51.715 70.68 51.885 ;
        RECT  1.14 48.915 70.68 49.085 ;
        RECT  1.14 46.115 70.68 46.285 ;
        RECT  1.14 43.315 70.68 43.485 ;
        RECT  1.14 40.515 70.68 40.685 ;
        RECT  1.14 37.715 70.68 37.885 ;
        RECT  1.14 34.915 70.68 35.085 ;
        RECT  1.14 32.115 70.68 32.285 ;
        RECT  1.14 29.315 70.68 29.485 ;
        RECT  1.14 26.515 70.68 26.685 ;
        RECT  1.14 23.715 70.68 23.885 ;
        RECT  1.14 20.915 70.68 21.085 ;
        RECT  1.14 18.115 70.68 18.285 ;
        RECT  1.14 15.315 70.68 15.485 ;
        RECT  1.14 12.515 70.68 12.685 ;
        RECT  1.14 9.715 70.68 9.885 ;
        RECT  1.14 6.915 70.68 7.085 ;
        RECT  1.14 4.115 70.68 4.285 ;
        RECT  1.14 1.315 70.68 1.485 ;
      VIA 59.14 203.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 203.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 203.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 203.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 203.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 203.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 163.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 123.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 83.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 208.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 208.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 208.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 205.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 205.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 205.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 203 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 203 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 203 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 200.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 200.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 200.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 197.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 197.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 197.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 194.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 194.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 194.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 191.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 191.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 191.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 189 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 189 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 189 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 186.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 186.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 186.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 183.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 183.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 183.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 180.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 180.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 180.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 177.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 177.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 177.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 175 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 175 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 175 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 172.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 172.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 172.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 208.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 208.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 208.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 205.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 205.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 205.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 203 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 203 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 203 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 200.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 200.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 200.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 197.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 197.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 197.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 194.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 194.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 194.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 191.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 191.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 191.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 189 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 189 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 189 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 186.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 186.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 186.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 183.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 183.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 183.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 180.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 180.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 180.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 177.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 177.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 177.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 175 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 175 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 175 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 172.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 172.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 172.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 169.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 169.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 166.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 166.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 163.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 163.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 161 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 161 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 161 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 158.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 158.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 155.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 155.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 152.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 152.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 149.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 149.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 147 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 147 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 147 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 144.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 144.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 141.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 141.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 138.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 138.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 135.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 135.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 133 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 133 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 133 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 130.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 130.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 127.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 127.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 124.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 124.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 121.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 121.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 119 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 119 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 119 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 116.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 116.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 113.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 113.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 110.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 110.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 107.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 107.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 105 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 105 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 105 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 102.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 102.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 99.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 99.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 96.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 96.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 93.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 93.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 91 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 91 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 91 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 88.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 88.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 85.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 85.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 82.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 82.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 79.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 79.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 77 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 77 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 77 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 74.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 74.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 71.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 71.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 68.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 68.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  30.9 2.715 31.38 210.085 ;
      LAYER metal1 ;
        RECT  1.14 209.915 70.68 210.085 ;
        RECT  1.14 207.115 70.68 207.285 ;
        RECT  1.14 204.315 70.68 204.485 ;
        RECT  1.14 201.515 70.68 201.685 ;
        RECT  1.14 198.715 70.68 198.885 ;
        RECT  1.14 195.915 70.68 196.085 ;
        RECT  1.14 193.115 70.68 193.285 ;
        RECT  1.14 190.315 70.68 190.485 ;
        RECT  1.14 187.515 70.68 187.685 ;
        RECT  1.14 184.715 70.68 184.885 ;
        RECT  1.14 181.915 70.68 182.085 ;
        RECT  1.14 179.115 70.68 179.285 ;
        RECT  1.14 176.315 70.68 176.485 ;
        RECT  1.14 173.515 70.68 173.685 ;
        RECT  1.14 170.715 70.68 170.885 ;
        RECT  1.14 167.915 70.68 168.085 ;
        RECT  1.14 165.115 70.68 165.285 ;
        RECT  1.14 162.315 70.68 162.485 ;
        RECT  1.14 159.515 70.68 159.685 ;
        RECT  1.14 156.715 70.68 156.885 ;
        RECT  1.14 153.915 70.68 154.085 ;
        RECT  1.14 151.115 70.68 151.285 ;
        RECT  1.14 148.315 70.68 148.485 ;
        RECT  1.14 145.515 70.68 145.685 ;
        RECT  1.14 142.715 70.68 142.885 ;
        RECT  1.14 139.915 70.68 140.085 ;
        RECT  1.14 137.115 70.68 137.285 ;
        RECT  1.14 134.315 70.68 134.485 ;
        RECT  1.14 131.515 70.68 131.685 ;
        RECT  1.14 128.715 70.68 128.885 ;
        RECT  1.14 125.915 70.68 126.085 ;
        RECT  1.14 123.115 70.68 123.285 ;
        RECT  1.14 120.315 70.68 120.485 ;
        RECT  1.14 117.515 70.68 117.685 ;
        RECT  1.14 114.715 70.68 114.885 ;
        RECT  1.14 111.915 70.68 112.085 ;
        RECT  1.14 109.115 70.68 109.285 ;
        RECT  1.14 106.315 70.68 106.485 ;
        RECT  1.14 103.515 70.68 103.685 ;
        RECT  1.14 100.715 70.68 100.885 ;
        RECT  1.14 97.915 70.68 98.085 ;
        RECT  1.14 95.115 70.68 95.285 ;
        RECT  1.14 92.315 70.68 92.485 ;
        RECT  1.14 89.515 70.68 89.685 ;
        RECT  1.14 86.715 70.68 86.885 ;
        RECT  1.14 83.915 70.68 84.085 ;
        RECT  1.14 81.115 70.68 81.285 ;
        RECT  1.14 78.315 70.68 78.485 ;
        RECT  1.14 75.515 70.68 75.685 ;
        RECT  1.14 72.715 70.68 72.885 ;
        RECT  1.14 69.915 70.68 70.085 ;
        RECT  1.14 67.115 70.68 67.285 ;
        RECT  1.14 64.315 70.68 64.485 ;
        RECT  1.14 61.515 70.68 61.685 ;
        RECT  1.14 58.715 70.68 58.885 ;
        RECT  1.14 55.915 70.68 56.085 ;
        RECT  1.14 53.115 70.68 53.285 ;
        RECT  1.14 50.315 70.68 50.485 ;
        RECT  1.14 47.515 70.68 47.685 ;
        RECT  1.14 44.715 70.68 44.885 ;
        RECT  1.14 41.915 70.68 42.085 ;
        RECT  1.14 39.115 70.68 39.285 ;
        RECT  1.14 36.315 70.68 36.485 ;
        RECT  1.14 33.515 70.68 33.685 ;
        RECT  1.14 30.715 70.68 30.885 ;
        RECT  1.14 27.915 70.68 28.085 ;
        RECT  1.14 25.115 70.68 25.285 ;
        RECT  1.14 22.315 70.68 22.485 ;
        RECT  1.14 19.515 70.68 19.685 ;
        RECT  1.14 16.715 70.68 16.885 ;
        RECT  1.14 13.915 70.68 14.085 ;
        RECT  1.14 11.115 70.68 11.285 ;
        RECT  1.14 8.315 70.68 8.485 ;
        RECT  1.14 5.515 70.68 5.685 ;
        RECT  1.14 2.715 70.68 2.885 ;
      VIA 31.14 210 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 210 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 210 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 207.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 207.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 207.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 204.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 204.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 204.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 201.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 201.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 201.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 198.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 198.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 198.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 196 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 196 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 196 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 193.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 193.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 193.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 190.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 190.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 190.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 187.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 187.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 187.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 184.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 184.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 184.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 182 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 182 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 182 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 179.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 179.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 179.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 176.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 176.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 176.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 173.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 173.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 173.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 170.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 170.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 170.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 168 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 168 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 168 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 165.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 165.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 162.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 162.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 159.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 159.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 156.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 156.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 154 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 154 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 154 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 151.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 151.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 148.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 148.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 145.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 145.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 142.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 142.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 140 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 140 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 140 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 137.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 137.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 134.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 134.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 131.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 131.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 128.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 128.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 126 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 126 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 126 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 123.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 123.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 120.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 120.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 117.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 117.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 114.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 114.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 112 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 112 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 112 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 109.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 109.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 106.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 106.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 103.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 103.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 100.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 100.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 98 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 98 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 98 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 95.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 95.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 92.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 92.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 89.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 89.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 86.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 86.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 84 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 84 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 84 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 81.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 81.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 78.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 78.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 75.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 75.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 72.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 72.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 70 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 70 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 70 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 169.68 0.14 169.82 ;
    END
  END clk
  PIN enable_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 95.2 0.14 95.34 ;
    END
  END enable_write
  PIN read_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 113.68 0.14 113.82 ;
    END
  END read_data[0]
  PIN read_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 106.4 71.785 106.54 ;
    END
  END read_data[1]
  PIN read_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 108.08 71.785 108.22 ;
    END
  END read_data[2]
  PIN read_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 108.64 71.785 108.78 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 112.56 0.14 112.7 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 113.68 71.785 113.82 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 113.12 71.785 113.26 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 107.52 71.785 107.66 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 106.96 71.785 107.1 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 113.12 0.14 113.26 ;
    END
  END read_data[9]
  PIN read_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 44.24 71.785 44.38 ;
    END
  END read_index[0]
  PIN read_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 45.36 71.785 45.5 ;
    END
  END read_index[1]
  PIN read_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 47.04 71.785 47.18 ;
    END
  END read_index[2]
  PIN read_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 94.64 0.14 94.78 ;
    END
  END read_index[3]
  PIN read_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 112 0.14 112.14 ;
    END
  END read_index[4]
  PIN read_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 112.56 71.785 112.7 ;
    END
  END read_index[5]
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 117.6 0.14 117.74 ;
    END
  END write_data[0]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 117.04 0.14 117.18 ;
    END
  END write_data[1]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 114.24 71.785 114.38 ;
    END
  END write_data[2]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 95.2 71.785 95.34 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 114.24 0.14 114.38 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 120.96 71.785 121.1 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 93.52 71.785 93.66 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 116.48 0.14 116.62 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 102.48 71.785 102.62 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  71.645 90.16 71.785 90.3 ;
    END
  END write_data[9]
  PIN write_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 95.76 0.14 95.9 ;
    END
  END write_index[0]
  PIN write_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 98 0.14 98.14 ;
    END
  END write_index[1]
  PIN write_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 97.44 0.14 97.58 ;
    END
  END write_index[2]
  PIN write_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 96.32 0.14 96.46 ;
    END
  END write_index[3]
  PIN write_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 96.88 0.14 97.02 ;
    END
  END write_index[4]
  PIN write_index[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 98.56 0.14 98.7 ;
    END
  END write_index[5]
  OBS
    LAYER metal1 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal2 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal3 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal4 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal5 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal6 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal7 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal8 ;
     RECT  0 1.315 71.785 210.085 ;
    LAYER metal9 ;
     RECT  0 1.315 71.785 210.085 ;
  END
END SmallBuffer64
END LIBRARY
