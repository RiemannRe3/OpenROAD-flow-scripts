VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO SmallBuffer32
  FOREIGN SmallBuffer32 0 0 ;
  CLASS BLOCK ;
  SIZE 113.645 BY 68.985 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 42.7 59.38 44.1 ;
        RECT  2.9 2.7 59.38 4.1 ;
      LAYER metal4 ;
        RECT  58.9 1.315 59.38 65.885 ;
        RECT  2.9 1.315 3.38 65.885 ;
      LAYER metal1 ;
        RECT  1.14 65.715 112.48 65.885 ;
        RECT  1.14 62.915 112.48 63.085 ;
        RECT  1.14 60.115 112.48 60.285 ;
        RECT  1.14 57.315 112.48 57.485 ;
        RECT  1.14 54.515 112.48 54.685 ;
        RECT  1.14 51.715 112.48 51.885 ;
        RECT  1.14 48.915 112.48 49.085 ;
        RECT  1.14 46.115 112.48 46.285 ;
        RECT  1.14 43.315 112.48 43.485 ;
        RECT  1.14 40.515 112.48 40.685 ;
        RECT  1.14 37.715 112.48 37.885 ;
        RECT  1.14 34.915 112.48 35.085 ;
        RECT  1.14 32.115 112.48 32.285 ;
        RECT  1.14 29.315 112.48 29.485 ;
        RECT  1.14 26.515 112.48 26.685 ;
        RECT  1.14 23.715 112.48 23.885 ;
        RECT  1.14 20.915 112.48 21.085 ;
        RECT  1.14 18.115 112.48 18.285 ;
        RECT  1.14 15.315 112.48 15.485 ;
        RECT  1.14 12.515 112.48 12.685 ;
        RECT  1.14 9.715 112.48 9.885 ;
        RECT  1.14 6.915 112.48 7.085 ;
        RECT  1.14 4.115 112.48 4.285 ;
        RECT  1.14 1.315 112.48 1.485 ;
      VIA 59.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.9 62.7 87.38 64.1 ;
        RECT  30.9 22.7 87.38 24.1 ;
      LAYER metal4 ;
        RECT  86.9 2.715 87.38 67.285 ;
        RECT  30.9 2.715 31.38 67.285 ;
      LAYER metal1 ;
        RECT  1.14 67.115 112.48 67.285 ;
        RECT  1.14 64.315 112.48 64.485 ;
        RECT  1.14 61.515 112.48 61.685 ;
        RECT  1.14 58.715 112.48 58.885 ;
        RECT  1.14 55.915 112.48 56.085 ;
        RECT  1.14 53.115 112.48 53.285 ;
        RECT  1.14 50.315 112.48 50.485 ;
        RECT  1.14 47.515 112.48 47.685 ;
        RECT  1.14 44.715 112.48 44.885 ;
        RECT  1.14 41.915 112.48 42.085 ;
        RECT  1.14 39.115 112.48 39.285 ;
        RECT  1.14 36.315 112.48 36.485 ;
        RECT  1.14 33.515 112.48 33.685 ;
        RECT  1.14 30.715 112.48 30.885 ;
        RECT  1.14 27.915 112.48 28.085 ;
        RECT  1.14 25.115 112.48 25.285 ;
        RECT  1.14 22.315 112.48 22.485 ;
        RECT  1.14 19.515 112.48 19.685 ;
        RECT  1.14 16.715 112.48 16.885 ;
        RECT  1.14 13.915 112.48 14.085 ;
        RECT  1.14 11.115 112.48 11.285 ;
        RECT  1.14 8.315 112.48 8.485 ;
        RECT  1.14 5.515 112.48 5.685 ;
        RECT  1.14 2.715 112.48 2.885 ;
      VIA 87.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 87.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 63.4 via4_5_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via6_7_960_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_960_2800_5_2_600_600 ;
      VIA 31.14 23.4 via4_5_960_2800_5_2_600_600 ;
      VIA 87.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 87.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 87.14 2.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 67.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 67.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 17.92 113.645 18.06 ;
    END
  END clk
  PIN enable_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  65.545 0 65.685 0.14 ;
    END
  END enable_write
  PIN read_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END read_data[0]
  PIN read_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END read_data[1]
  PIN read_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.105 0 66.245 0.14 ;
    END
  END read_data[2]
  PIN read_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  64.985 68.845 65.125 68.985 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  58.825 68.845 58.965 68.985 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  56.025 68.845 56.165 68.985 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  65.545 68.845 65.685 68.985 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  62.745 68.845 62.885 68.985 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  57.145 0 57.285 0.14 ;
    END
  END read_data[9]
  PIN read_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 19.04 113.645 19.18 ;
    END
  END read_index[0]
  PIN read_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 20.16 113.645 20.3 ;
    END
  END read_index[1]
  PIN read_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 23.52 113.645 23.66 ;
    END
  END read_index[2]
  PIN read_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 45.36 0.14 45.5 ;
    END
  END read_index[3]
  PIN read_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  62.185 68.845 62.325 68.985 ;
    END
  END read_index[4]
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 41.44 0.14 41.58 ;
    END
  END write_data[0]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 30.8 113.645 30.94 ;
    END
  END write_data[1]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 48.16 0.14 48.3 ;
    END
  END write_data[2]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 38.08 0.14 38.22 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 32.48 113.645 32.62 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 44.24 0.14 44.38 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 46.48 0.14 46.62 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 26.88 113.645 27.02 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 42 0.14 42.14 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  113.505 28 113.645 28.14 ;
    END
  END write_data[9]
  PIN write_index[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  67.225 0 67.365 0.14 ;
    END
  END write_index[0]
  PIN write_index[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END write_index[1]
  PIN write_index[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END write_index[2]
  PIN write_index[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END write_index[3]
  PIN write_index[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.305 0 49.445 0.14 ;
    END
  END write_index[4]
  OBS
    LAYER metal1 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal2 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal3 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal4 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal5 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal6 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal7 ;
     RECT  0 0 113.645 68.985 ;
    LAYER metal9 ;
     RECT  0 0 113.645 68.985 ;
  END
END SmallBuffer32
END LIBRARY
